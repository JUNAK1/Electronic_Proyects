LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.numeric_std.all;

ENTITY ROM IS
	generic (
		DATA_WIDTH : natural := 15;--19
		ADDR_WIDTH : natural := 4--3
);
	PORT (
		clock: IN STD_LOGIC;
		data: OUT STD_LOGIC_VECTOR (DATA_WIDTH-1 DOWNTO 0);
		add: IN STD_LOGIC_VECTOR(ADDR_WIDTH-1 DOWNTO 0)
	);
END ROM;

ARCHITECTURE rtl OF ROM IS
	SUBTYPE datos IS STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0);
	TYPE rom_type IS ARRAY(0 to (2**ADDR_WIDTH)-1) OF datos;
	SIGNAL ROM: ROM_TYPE :=(		
"010000000100000","101000000000101","010000001011000","110100000000101",
"101000000001010","110000000000101","110110000001010","101000000001111",
"010000110010000","110010000000000","000000000000000","000000000000000",
"000000000000000","000000000000000","000000000000000","000000000000000");	
BEGIN
	PROCESS (clock)
	BEGIN
		IF (RISING_EDGE(clock)) THEN	
			data <= ROM(conv_integer(add));
		END IF;
	END PROCESS;

END rtl;